LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY Decoder IS
	PORT (
		OPCODE : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		FUNCT : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		OPERACAO : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		OUTPUT : OUT STD_LOGIC_VECTOR(10 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE arch_name OF Decoder IS
	CONSTANT ADDR : STD_LOGIC_VECTOR(5 DOWNTO 0) := "100000";
	CONSTANT SUBR : STD_LOGIC_VECTOR(5 DOWNTO 0) := "100111";
	CONSTANT LW : STD_LOGIC_VECTOR(5 DOWNTO 0) := "100011";
	CONSTANT SW : STD_LOGIC_VECTOR(5 DOWNTO 0) := "101011";
	CONSTANT BEQ : STD_LOGIC_VECTOR(5 DOWNTO 0) := "000100";
	CONSTANT J : STD_LOGIC_VECTOR(5 DOWNTO 0) := "000010";
	-- TipoR|SelMuxJump|SelMuxRtRd|write_REG(1)|habMUX(rt/imediato)|OP(2)|SelMuxMEMULA|habFlagEqual|
	--read_RAM|write_RAM
BEGIN

	OUTPUT <= "0" & "0011" & OPERACAO & "1010" WHEN (OPCODE = LW) ELSE
		"0" & "0001"  & OPERACAO & "1001" WHEN (OPCODE = SW) ELSE
		"0" & "0000" & OPERACAO & "1100" WHEN (OPCODE = BEQ) ELSE
		"1" & "0110" & OPERACAO & "0000" WHEN (FUNCT = ADDR AND OPCODE = "000000") ELSE
		"1" & "0110" & OPERACAO & "0000" WHEN (FUNCT = SUBR AND OPCODE = "000000") ELSE
		"0" & "1000" & OPERACAO & "0000" WHEN (OPCODE = J) ELSE
		"00000000000";
END ARCHITECTURE;