LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY Decoder IS
	PORT (
		OPCODE : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		FUNCT : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		OPERACAO : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		OUTPUT : OUT STD_LOGIC_VECTOR(13 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE arch_name OF Decoder IS
	CONSTANT ADDR : STD_LOGIC_VECTOR(5 DOWNTO 0) := "100000";
	CONSTANT SUBR : STD_LOGIC_VECTOR(5 DOWNTO 0) := "100010";
	CONSTANT LW : STD_LOGIC_VECTOR(5 DOWNTO 0) := "100011";
	CONSTANT SW : STD_LOGIC_VECTOR(5 DOWNTO 0) := "101011";
	CONSTANT BEQ : STD_LOGIC_VECTOR(5 DOWNTO 0) := "000100";
	CONSTANT J : STD_LOGIC_VECTOR(5 DOWNTO 0) := "000010";
	CONSTANT SLT : STD_LOGIC_VECTOR(5 DOWNTO 0) := "101010";
	CONSTANT ANDR : STD_LOGIC_VECTOR(5 DOWNTO 0) := "100100";
	CONSTANT ORR : STD_LOGIC_VECTOR(5 DOWNTO 0) := "100101";

	CONSTANT ORI : STD_LOGIC_VECTOR(5 DOWNTO 0) := "001101";
	CONSTANT ADDI : STD_LOGIC_VECTOR(5 DOWNTO 0) := "001000";
	CONSTANT ANDI : STD_LOGIC_VECTOR(5 DOWNTO 0) := "001100";
	CONSTANT SLTI : STD_LOGIC_VECTOR(5 DOWNTO 0) := "001010";
	
	CONSTANT JAL : STD_LOGIC_VECTOR(5 DOWNTO 0) := "000011";
	CONSTANT JR : STD_LOGIC_VECTOR(5 DOWNTO 0) := "001000";
	CONSTANT LUI : STD_LOGIC_VECTOR(5 DOWNTO 0) := "001111";
	CONSTANT BNE : STD_LOGIC_VECTOR(5 DOWNTO 0) := "000101";

-- JR|SelMuxBEQJmp|muxRTRD|ORI_ANDI|habEscritaReg|muxRTImediato|TipoR|muxULAMEM|BEQ|BNE|Leitura|Escrita
BEGIN

	OUTPUT <= "0" & "000011" & "0" & "01" & "0010" WHEN (OPCODE = LW) ELSE
			  "0" & "000001" & "0" & "00" & "0001" WHEN (OPCODE = SW) ELSE
			  "0" & "000000" & "0" & "00" & "1000" WHEN (OPCODE = BEQ) ELSE
			  "0" & "000000" & "0" & "00" & "0100" WHEN (OPCODE = BNE) ELSE
			  "0" & "001010" & "1" & "00" & "0000" WHEN (((FUNCT = ADDR) OR (FUNCT = SUBR) OR (FUNCT = ORR) OR (FUNCT = ANDR) OR (FUNCT = SLT)) AND OPCODE = "000000") ELSE 
			  "0" & "000011" & "0" & "00" & "0000" WHEN ((OPCODE = ADDI) OR (OPCODE = SLTI)) ELSE
			  "0" & "000111" & "0" & "00" & "0000" WHEN ((OPCODE = ORI) OR (OPCODE = ANDI)) ELSE
			  "0" & "100000" & "0" & "00" & "0000" WHEN (OPCODE = J) ELSE
			  "0" & "000010" & "0" & "11" & "0000" WHEN (OPCODE = LUI) ELSE
			  "0" & "110010" & "0" & "10" & "0000" WHEN (OPCODE = JAL) ELSE
			  "1" & "000000" & "1" & "00" & "0000" WHEN (FUNCT = JR) ELSE
			  ---- FALTA ESCREVER OS DECODERS DO JAL, JR E IR NO DECODER OPCODE E DEBUG MONITOR MUDAR O MUXRTRD
			  "00000000000000";
END ARCHITECTURE;