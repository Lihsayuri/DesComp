library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 15;
          addrWidth: natural := 9
    );
   port (
          Endereco : in std_logic_vector (8 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI : std_logic_vector(3 downto 0) := "0100";
  constant STA : std_logic_vector(3 downto 0) := "0101";
  constant JMP : std_logic_vector(3 downto 0) := "0110";
  constant JEQ : std_logic_vector(3 downto 0) := "0111";
  constant CEQ : std_logic_vector(3 downto 0) := "1000";
  constant JSR : std_logic_vector(3 downto 0) := "1001";
  constant RET : std_logic_vector(3 downto 0) := "1010";
  constant ANDI : std_logic_vector(3 downto 0) := "1011";
  constant CLT : std_logic_vector (3 downto 0) := "1100"; -- CLT
  constant JLT : std_logic_vector (3 downto 0) := "1101"; -- JLT. OBS: ainda temos 1110 e 1111
  constant ADDI : std_logic_vector (3 downto 0) := "1110"; 
  constant SUBI : std_logic_vector (3 downto 0) := "1111";

  
  constant R0:    std_logic_vector (1 DOWNTO 0)	:= "00";
  constant R1:    std_logic_vector (1 DOWNTO 0)	:= "01";
  constant R2:    std_logic_vector (1 DOWNTO 0)	:= "10";
  constant R3:    std_logic_vector (1 DOWNTO 0)	:= "11";

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
		
  begin
      -- Palavra de Controle = SelMUX, Habilita_A, Reset_A, Operacao_ULA
					-- Inicializa os endereços:
					
						-- SETUP: INICIALIZAÇÃO DE ENDEREÇOS E ALGUMAS VARIÁVEIS
		tmp(0) := LDI  &  R0  &  '0'  &  x"00";	-- LDI $0, R0      	# Inicializando algumas variáveis importantes : R0 = 0
		tmp(1) := LDI  &  R1  &  '0'  &  x"01";	-- LDI $1, R1      	# R1 = 1
		tmp(2) := LDI  &  R2  &  '0'  &  x"06";	-- LDI $6, R2      	# R2 = 6
		tmp(3) := LDI  &  R3  &  '0'  &  x"0a";	-- LDI $10, R3     	# R3 = 10
		tmp(4) := STA  &  R0  &  '1'  &  x"00";	-- STA @256, R0    	# Armazena o valor do R0 no LEDR0 ~ LEDR7
		tmp(5) := STA  &  R0  &  '1'  &  x"01";	-- STA @257, R0    	# Armazena o valor do R0 no LEDR8
		tmp(6) := STA  &  R0  &  '1'  &  x"02";	-- STA @258, R0    	# Armazena o valor do R0 no LEDR9
		tmp(7) := STA  &  R0  &  '1'  &  x"20";	-- STA @288, R0    	# Armazena o valor do R0 no HEX0
		tmp(8) := STA  &  R0  &  '1'  &  x"21";	-- STA @289, R0    	# Armazena o valor do R0 no HEX1
		tmp(9) := STA  &  R0  &  '1'  &  x"22";	-- STA @290, R0    	# Armazena o valor do R0 no HEX2
		tmp(10) := STA  &  R0  &  '1'  &  x"23";	-- STA @291, R0    	# Armazena o valor do R0 no HEX3
		tmp(11) := STA  &  R0  &  '1'  &  x"24";	-- STA @292, R0    	# Armazena o valor do R0 no HEX4
		tmp(12) := STA  &  R0  &  '1'  &  x"25";	-- STA @293, R0    	# Armazena o valor do R0 no HEX5
		tmp(13) := STA  &  R0  &  '0'  &  x"00";	-- STA @0, R0      	# Armazena o valor do R0 em MEM[0] (unidades de segundo)
		tmp(14) := STA  &  R0  &  '0'  &  x"01";	-- STA @1, R0      	# Armazena o valor do R0 em MEM[1] (dezenas de segundo)
		tmp(15) := STA  &  R0  &  '0'  &  x"02";	-- STA @2, R0      	# Armazena o valor do R0 em MEM[2] (unidades de minuto)
		tmp(16) := STA  &  R0  &  '0'  &  x"03";	-- STA @3, R0      	# Armazena o valor do R0 em MEM[3] (dezenas de minuto)
		tmp(17) := STA  &  R0  &  '0'  &  x"04";	-- STA @4, R0      	# Armazena o valor do R0 em MEM[4] (unidades de hora)
		tmp(18) := STA  &  R0  &  '0'  &  x"05";	-- STA @5, R0      	# Armazena o valor do R0 em MEM[5] (dezenas de hora)
		tmp(19) := STA  &  R0  &  '0'  &  x"06";	-- STA @6, R0      	# Armazena o valor do R0 em MEM[6] (flag do despertador)
		tmp(20) := STA  &  R0  &  '0'  &  x"07";	-- STA @7, R0      	# Armazena o valor do R0 em MEM[7] (variável 0 para comparações)
		tmp(21) := STA  &  R1  &  '0'  &  x"08";	-- STA @8, R1      	# Armazena o valor do R1 em MEM[8] (variável 1 para incremento)
		tmp(22) := STA  &  R3  &  '0'  &  x"09";	-- STA @9, R3      	# Armazena o valor do R3 em MEM[9] (variável 10 para comparações)
		tmp(23) := STA  &  R2  &  '0'  &  x"0a";	-- STA @10, R2     	# Armazena o valor do R2 em MEM[10] (valor do despertador para UNIDADE DE SEGUNDO)
		tmp(24) := STA  &  R2  &  '0'  &  x"0b";	-- STA @11, R2     	# Armazena o valor do R2 em MEM[11] (valor do despertador para DEZENA DE SEGUNDO)
		tmp(25) := STA  &  R2  &  '0'  &  x"0c";	-- STA @12, R2     	# Armazena o valor do R2 em MEM[12] (valor do despertador para UNIDADE DE MINUTO)
		tmp(26) := STA  &  R2  &  '0'  &  x"0d";	-- STA @13, R2     	# Armazena o valor do R2 em MEM[13] (valor do despertador para DEZENA DE MINUTO)
		tmp(27) := STA  &  R2  &  '0'  &  x"0e";	-- STA @14, R2     	# Armazena o valor do R2 em MEM[14] (valor do despertador para UNIDADE DE HORA)
		tmp(28) := STA  &  R2  &  '0'  &  x"0f";	-- STA @15, R2     	# Armazena o valor do R2 em MEM[15] (valor do despertador para DEZENA DE HORA)
		tmp(29) := STA  &  R2  &  '0'  &  x"10";	-- STA @16, R2     	# Armazena o valor do R2 em MEM[16] (constante 6)
		tmp(30) := LDI  &  R0  &  '0'  &  x"02";	-- LDI $2, R0      	# Carrega 2 no registrador R0
		tmp(31) := STA  &  R0  &  '0'  &  x"11";	-- STA @17, R0     	# Armazena o valor do R0 em MEM[17] (constante 2)
		tmp(32) := LDI  &  R0  &  '0'  &  x"04";	-- LDI $4, R0      	# Carrega 4 no registrador R0
		tmp(33) := STA  &  R0  &  '0'  &  x"12";	-- STA @18, R0     	# Armazena o valor do R0 em MEM[18] (constante 4)
		tmp(34) := LDI  &  R0  &  '0'  &  x"18";	-- LDI $24, R0     	# Carrega 24 no registrador R0
		tmp(35) := STA  &  R0  &  '0'  &  x"13";	-- STA @19, R0     	# Armazena o valor do R0 em MEM[19] (constante 24)
		tmp(36) := NOP  &  R0  &  '0'  &  x"00";	-- NOP              	# LOOP PRINCIPAL
		tmp(37) := LDA  &  R0  &  '1'  &  x"60";	-- LDA @352, R0     	# Carrega o R0 com a leitura do botão KEY0
		tmp(38) := ANDI  &  R0  &  '0'  &  x"01";	-- ANDI @1, R0      	# Aplica máscara na leitura do botão
		tmp(39) := CEQ  &  R0  &  '0'  &  x"07";	-- CEQ @7, R0       	# Compara com 0
		tmp(40) := JEQ  &  R0  &  '0'  &  x"2b";	-- JEQ @LEITURA_KEY1 	# Se for 0, vai ler a próxima chave
		tmp(41) := JSR  &  R0  &  '0'  &  x"45";	-- JSR @INCREMENTO  	# Se for 1, vai pra sub-rotina de incremento
		tmp(42) := NOP  &  R0  &  '0'  &  x"00";	-- NOP              	# Aqui é onde o RET volta
		tmp(43) := LDA  &  R1  &  '1'  &  x"61";	-- LDA @353, R1     	# Carrega o R1 com a leitura do botão KEY1
		tmp(44) := ANDI  &  R1  &  '0'  &  x"01";	-- ANDI @1, R1      	# Aplica máscara na leitura do botão
		tmp(45) := CEQ  &  R1  &  '0'  &  x"07";	-- CEQ @7, R1       	# Compara com 0
		tmp(46) := JEQ  &  R0  &  '0'  &  x"31";	-- JEQ @CHAMA_CONFERE_LIMITE 	# Se for 0, vai conferir o limite 
		tmp(47) := JSR  &  R0  &  '0'  &  x"bb";	-- JSR @CONFIG_DESPERTADOR   	# Se for 1, vai pra sub-rotina de configuração do despertador
		tmp(48) := NOP  &  R0  &  '0'  &  x"00";	-- NOP              	# Aqui é onde o RET volta
		tmp(49) := JSR  &  R0  &  '0'  &  x"a0";	-- JSR @CONFERE_LIMITE  	# Chama a sub-rotina para verificar o limite
		tmp(50) := NOP  &  R0  &  '0'  &  x"00";	-- NOP              	# Aqui é onde o RET volta
		tmp(51) := LDA  &  R0  &  '1'  &  x"62";	-- LDA @354, R0    	# Carrega R2 com a leitura de KEY2
		tmp(52) := ANDI  &  R0  &  '0'  &  x"01";	-- ANDI @1, R0     	# Depois de fazer a leitura do botão aplica a máscara
		tmp(53) := CEQ  &  R0  &  '0'  &  x"07";	-- CEQ @7, R0      	# Compara com 0
		tmp(54) := JEQ  &  R0  &  '0'  &  x"38";	-- JEQ @LEITURA_KEY3 	# Se for 0, vai ler a próxima chave 
		tmp(55) := JSR  &  R0  &  '1'  &  x"28";	-- JSR @DESLIGA_DESPERTADOR 	# Se for 1, vai para a sub-rotina de configurar hora
		tmp(56) := LDA  &  R2  &  '1'  &  x"63";	-- LDA @355, R2    	# Carrega R2 com a leitura de KEY3
		tmp(57) := ANDI  &  R2  &  '0'  &  x"01";	-- ANDI @1, R2     	# Depois de fazer a leitura do botão aplica a máscara
		tmp(58) := CEQ  &  R2  &  '0'  &  x"07";	-- CEQ @7, R2      	# Compara com 0
		tmp(59) := JEQ  &  R0  &  '0'  &  x"3e";	-- JEQ @LEITURA_RESET 	# Se for 0, vai ler a próxima chave 
		tmp(60) := JSR  &  R0  &  '1'  &  x"35";	-- JSR @CONFIGURA_HORARIO 	# Se for 1, vai para a sub-rotina de configurar hora
		tmp(61) := NOP  &  R0  &  '0'  &  x"00";	-- NOP
		tmp(62) := LDA  &  R3  &  '1'  &  x"64";	-- LDA @356, R3     	# Carrega o R3 com a leitura do botão FPGA_RESET 
		tmp(63) := ANDI  &  R3  &  '0'  &  x"01";	-- ANDI @1, R3      	# Aplica máscara na leitura do botão
		tmp(64) := CEQ  &  R3  &  '0'  &  x"08";	-- CEQ @8, R3       	# Compara com 1
		tmp(65) := JEQ  &  R0  &  '0'  &  x"43";	-- JEQ @CHAMA_ATUALIZA_DISPLAY 	# Se for 1, vai pra subrotina pra reiniciar a contagem (botão é o contrário. 0 - ativado. 1 - desativado)
		tmp(66) := JSR  &  R0  &  '0'  &  x"95";	-- JSR @REINICIAR_CONTAGEM  	# Chama sub-rotina de reiniciar a contagem
		tmp(67) := JSR  &  R0  &  '0'  &  x"83";	-- JSR @ATUALIZA_SEVEN_SEG  	# Chama sub-rotina de atualizar o display de sete segmentos
		tmp(68) := JMP  &  R0  &  '0'  &  x"24";	-- JMP @LOOP_PRINCIPAL      	# Volta para o início do loop principal
		tmp(69) := STA  &  R0  &  '1'  &  x"ff";	-- STA @511, R0     	# Limpa a leitura do botão KEY0
		tmp(70) := LDA  &  R0  &  '0'  &  x"00";	-- LDA @0, R0       	# Carrega o valor das unidades de segundo em R0
		tmp(71) := ADDI  &  R0  &  '0'  &  x"01";	-- ADDI $1, R0      	# Soma com 1 e guarda resultado em R0
		tmp(72) := CEQ  &  R0  &  '0'  &  x"09";	-- CEQ @9, R0       	# Compara com 10
		tmp(73) := JEQ  &  R0  &  '0'  &  x"4c";	-- JEQ @INC_DEZENA  	# Se for 10, vai para as dezenas de segundo
		tmp(74) := STA  &  R0  &  '0'  &  x"00";	-- STA @0, R0       	# Se não, armazena o valor das unidades de segundo
		tmp(75) := JMP  &  R0  &  '0'  &  x"82";	-- JMP @FIM_INCREMENTO 	# E retorna
		tmp(76) := LDA  &  R0  &  '0'  &  x"07";	-- LDA @7, R0      	# Carrega 0 no R0
		tmp(77) := STA  &  R0  &  '0'  &  x"00";	-- STA @0, R0      	# Carrega 0 nas unidades de segundo
		tmp(78) := LDA  &  R0  &  '0'  &  x"01";	-- LDA @1, R0      	# Carrega o valor das dezenas de segundo em R0
		tmp(79) := ADDI  &  R0  &  '0'  &  x"01";	-- ADDI $1, R0     	# Soma com 1 e guarda resultado em R0
		tmp(80) := CEQ  &  R0  &  '0'  &  x"10";	-- CEQ @16, R0      	# Compara com 6
		tmp(81) := JEQ  &  R0  &  '0'  &  x"54";	-- JEQ @INC_CENTENA 	# Se for 6, vai para as unidades de minuto
		tmp(82) := STA  &  R0  &  '0'  &  x"01";	-- STA @1, R0      	# Se não, armazena o valor das dezenas de segundo
		tmp(83) := JMP  &  R0  &  '0'  &  x"82";	-- JMP @FIM_INCREMENTO 	# E retorna
		tmp(84) := LDA  &  R0  &  '0'  &  x"07";	-- LDA @7, R0      	# Carrega 0 no R0
		tmp(85) := STA  &  R0  &  '0'  &  x"01";	-- STA @1, R0      	# Carrega 0 nas dezenas de segundo
		tmp(86) := LDA  &  R0  &  '0'  &  x"02";	-- LDA @2, R0      	# Carrega o valor das unidades de minuto em R0
		tmp(87) := ADDI  &  R0  &  '0'  &  x"01";	-- ADDI $1, R0     	# Soma com 1 e guarda resultado em R0
		tmp(88) := CEQ  &  R0  &  '0'  &  x"09";	-- CEQ @9, R0      	# Compara com 10
		tmp(89) := JEQ  &  R0  &  '0'  &  x"5c";	-- JEQ @INC_MILHAR 	# Se for 10, vai para as dezenas de minuto
		tmp(90) := STA  &  R0  &  '0'  &  x"02";	-- STA @2, R0      	# Se não, armazena o valor das unidades de minuto
		tmp(91) := JMP  &  R0  &  '0'  &  x"82";	-- JMP @FIM_INCREMENTO 	# E retorna
		tmp(92) := LDA  &  R0  &  '0'  &  x"07";	-- LDA @7, R0      	# Carrega 0 no R0
		tmp(93) := STA  &  R0  &  '0'  &  x"02";	-- STA @2, R0      	# Carrega 0 nas unidades de minuto
		tmp(94) := LDA  &  R0  &  '0'  &  x"03";	-- LDA @3, R0      	# Carrega o valor das dezenas de minuto em R0
		tmp(95) := ADDI  &  R0  &  '0'  &  x"01";	-- ADDI $1, R0     	# Soma com 1 e guarda resultado em R0
		tmp(96) := CEQ  &  R0  &  '0'  &  x"10";	-- CEQ @16, R0      	# Compara com 6
		tmp(97) := JEQ  &  R0  &  '0'  &  x"64";	-- JEQ @INC_DEZMILHAR  	# Se for 6, vai para as unidades de hora
		tmp(98) := STA  &  R0  &  '0'  &  x"03";	-- STA @3, R0      	# Se não, armazena o valor das dezenas de minuto
		tmp(99) := JMP  &  R0  &  '0'  &  x"82";	-- JMP @FIM_INCREMENTO 	# E retorna
		tmp(100) := LDA  &  R0  &  '0'  &  x"07";	-- LDA @7, R0      	# Carrega 0 no R0
		tmp(101) := STA  &  R0  &  '0'  &  x"03";	-- STA @3, R0      	# Carrega 0 nas dezenas de minuto
		tmp(102) := LDA  &  R0  &  '0'  &  x"04";	-- LDA @4, R0      	# Carrega o valor das unidades de hora
		tmp(103) := ADDI  &  R0  &  '0'  &  x"01";	-- ADDI $1, R0     	# Soma com 1 e guarda resultado em R0
		tmp(104) := CEQ  &  R0  &  '0'  &  x"12";	-- CEQ @18, R0     	# Compara com 4
		tmp(105) := JEQ  &  R0  &  '0'  &  x"6e";	-- JEQ @CONFERE_24 	# Se for 4, vai conferir se as dezenas de hora são 2
		tmp(106) := CEQ  &  R0  &  '0'  &  x"09";	-- CEQ @9, R0      	# Caso contrário compara com 10
		tmp(107) := JEQ  &  R0  &  '0'  &  x"75";	-- JEQ @INC_CENTMILHAR 	# Se for igual a 10, vai para as dezenas de hora
		tmp(108) := STA  &  R0  &  '0'  &  x"04";	-- STA @4, R0      	# Caso contrário, armazena o valor das unidades de hora
		tmp(109) := JMP  &  R0  &  '0'  &  x"82";	-- JMP @FIM_INCREMENTO 	# E retorna
		tmp(110) := LDA  &  R1  &  '0'  &  x"05";	-- LDA @5, R1      	#Carrega o valor das dezenas de hora
		tmp(111) := CEQ  &  R1  &  '0'  &  x"11";	-- CEQ @17, R1     	# Compara com 2
		tmp(112) := JEQ  &  R0  &  '0'  &  x"7b";	-- JEQ @REINICIAR_CONTAGEM_24 	# Se for 2, daí deu 24h de fato
		tmp(113) := CEQ  &  R0  &  '0'  &  x"09";	-- CEQ @9, R0      	# Caso contrário compara com 10
		tmp(114) := JEQ  &  R0  &  '0'  &  x"75";	-- JEQ @INC_CENTMILHAR 	# Se for igual a 10, vai para as dezenas de hora
		tmp(115) := STA  &  R0  &  '0'  &  x"04";	-- STA @4, R0      	# Caso contrário, armazena o valor das unidades de hora
		tmp(116) := JMP  &  R0  &  '0'  &  x"82";	-- JMP @FIM_INCREMENTO
		tmp(117) := LDA  &  R0  &  '0'  &  x"07";	-- LDA @7, R0      	# Carrega 0 no R0
		tmp(118) := STA  &  R0  &  '0'  &  x"04";	-- STA @4, R0      	# Carrega 0 nas unidades de hora 
		tmp(119) := LDA  &  R0  &  '0'  &  x"05";	-- LDA @5, R0      	# Carrega o valor das dezenas de hora
		tmp(120) := ADDI  &  R0  &  '0'  &  x"01";	-- ADDI $1, R0     	# Soma com 1 e guarda resultado em R0
		tmp(121) := STA  &  R0  &  '0'  &  x"05";	-- STA @5, R0      	# Armazena o valor das centena de milhar
		tmp(122) := JMP  &  R0  &  '0'  &  x"82";	-- JMP @FIM_INCREMENTO
		tmp(123) := LDA  &  R0  &  '0'  &  x"07";	-- LDA @7, R0      	# Carrega o R0 com o valor 0
		tmp(124) := STA  &  R0  &  '0'  &  x"00";	-- STA @0, R0      	#  Armazena o valor 0 nas unidades de segundo
		tmp(125) := STA  &  R0  &  '0'  &  x"01";	-- STA @1, R0      	#  Armazena o valor 0 nas dezenas
		tmp(126) := STA  &  R0  &  '0'  &  x"02";	-- STA @2, R0      	#  Armazena o valor 0 nas centenas
		tmp(127) := STA  &  R0  &  '0'  &  x"03";	-- STA @3, R0      	#  Armazena o valor 0 nos milhares
		tmp(128) := STA  &  R0  &  '0'  &  x"04";	-- STA @4, R0      	#  Armazena o valor 0 nas dezenas de milhar
		tmp(129) := STA  &  R0  &  '0'  &  x"05";	-- STA @5, R0      	#  Armazena o valor 0 nas centenas de milhar
		tmp(130) := RET  &  R0  &  '0'  &  x"00";	-- RET
		tmp(131) := LDA  &  R0  &  '0'  &  x"00";	-- LDA @0, R0      	# Carrega o valor das unidades de segundo em R0
		tmp(132) := LDA  &  R1  &  '0'  &  x"01";	-- LDA @1, R1      	# Carrega o valor das dezenas  de segundo em R1
		tmp(133) := LDA  &  R2  &  '0'  &  x"02";	-- LDA @2, R2      	# Carrega o valor das unidades de minuto em R2
		tmp(134) := STA  &  R0  &  '1'  &  x"20";	-- STA @288, R0    	# Guarda o valor das unidades de segundo no HEX0
		tmp(135) := STA  &  R1  &  '1'  &  x"21";	-- STA @289, R1    	# Guarda o valor das dezenas de segundo no HEX1 
		tmp(136) := STA  &  R2  &  '1'  &  x"22";	-- STA @290, R2    	# Guarda o valor das unidades de minuto no HEX2
		tmp(137) := LDA  &  R0  &  '0'  &  x"03";	-- LDA @3, R0      	# Carrega o valor das dezenas de minuto em R0
		tmp(138) := LDA  &  R1  &  '0'  &  x"04";	-- LDA @4, R1      	# Carrega o valor das unidades de hora em R1
		tmp(139) := LDA  &  R2  &  '0'  &  x"05";	-- LDA @5, R2      	# Carrega o valor das dezenas de hora em R2
		tmp(140) := STA  &  R0  &  '1'  &  x"23";	-- STA @291, R0    	# Guarda o valor das dezenas de minuto no HEX3
		tmp(141) := STA  &  R1  &  '1'  &  x"24";	-- STA @292, R1    	# Guarda o valor das unidades de hora no HEX4
		tmp(142) := STA  &  R2  &  '1'  &  x"25";	-- STA @293, R2    	# Guarda o valor das dezenas de hora no HEX5
		tmp(143) := LDA  &  R0  &  '0'  &  x"06";	-- LDA @6, R0      	# Carrega o valor da flag do despertador 
		tmp(144) := CEQ  &  R0  &  '0'  &  x"07";	-- CEQ @7, R0      	# Compara o valor da flag com 0
		tmp(145) := JEQ  &  R0  &  '0'  &  x"94";	-- JEQ @FIM_ATUALIZA_TELA 	# Se for 0 a flag está inativa: então termina sub-rotina
		tmp(146) := LDA  &  R2  &  '0'  &  x"08";	-- LDA @8, R2      	# Caso contrário, carrega 1 em R2
		tmp(147) := STA  &  R2  &  '1'  &  x"01";	-- STA @257, R2    	# Salva o 1 no LEDR8
		tmp(148) := RET  &  R0  &  '0'  &  x"00";	-- RET
		tmp(149) := LDA  &  R0  &  '0'  &  x"07";	-- LDA @7, R0      	# Carrega o R0 com o valor 0
		tmp(150) := STA  &  R0  &  '0'  &  x"00";	-- STA @0, R0      	# Armazena o valor 0 nas unidades de segundo
		tmp(151) := STA  &  R0  &  '0'  &  x"01";	-- STA @1, R0      	# Armazena o valor 0 nas dezenas de segundo
		tmp(152) := STA  &  R0  &  '0'  &  x"02";	-- STA @2, R0      	# Armazena o valor 0 nas unidades de minuto
		tmp(153) := STA  &  R0  &  '0'  &  x"03";	-- STA @3, R0      	# Armazena o valor 0 nas dezenas de minuto
		tmp(154) := STA  &  R0  &  '0'  &  x"04";	-- STA @4, R0      	# Armazena o valor 0 nas unidades de hora
		tmp(155) := STA  &  R0  &  '0'  &  x"05";	-- STA @5, R0      	# Armazena o valor 0 nas dezenas de hora
		tmp(156) := STA  &  R0  &  '0'  &  x"06";	-- STA @6, R0      	# Armazena o valor 0 na flag do despertador
		tmp(157) := STA  &  R0  &  '1'  &  x"01";	-- STA @257, R0    	# Armazena o valor 0 no LEDR8
		tmp(158) := STA  &  R0  &  '1'  &  x"02";	-- STA @258, R0    	# Armazena o valor 0 no LEDR9
		tmp(159) := RET  &  R0  &  '0'  &  x"00";	-- RET
		tmp(160) := LDA  &  R0  &  '0'  &  x"0a";	-- LDA @10, R0      	# Carrega o valor do limite das unidades de segundo em R0
		tmp(161) := CEQ  &  R0  &  '0'  &  x"00";	-- CEQ @0, R0     	# Compara com as unidades de segundo
		tmp(162) := JEQ  &  R0  &  '0'  &  x"a4";	-- JEQ @CONFERE_LIMITE_SEG2 	# Se for igual, vai conferir as dezenas de segundo
		tmp(163) := JMP  &  R0  &  '0'  &  x"ba";	-- JMP @FIM_CONFERE_LIMITE   	# Caso o contrário já retorna
		tmp(164) := LDA  &  R1  &  '0'  &  x"0b";	-- LDA @11, R1      	# Carrega o valor do limite das dezenas de segundo em R1
		tmp(165) := CEQ  &  R1  &  '0'  &  x"01";	-- CEQ @1, R1     	# Compara com as dezenas de segundo
		tmp(166) := JEQ  &  R0  &  '0'  &  x"a8";	-- JEQ @CONFERE_LIMITE_MIN1 	# Se for igual, vai conferir as unidades de minuto
		tmp(167) := JMP  &  R0  &  '0'  &  x"ba";	-- JMP @FIM_CONFERE_LIMITE   	# Caso o contrário já retorna
		tmp(168) := LDA  &  R2  &  '0'  &  x"0c";	-- LDA @12, R2      	# Carrega o valor do limite das unidades de minuto em R2
		tmp(169) := CEQ  &  R2  &  '0'  &  x"02";	-- CEQ @2, R2     	# Compara com as unidades de minuto
		tmp(170) := JEQ  &  R0  &  '0'  &  x"ac";	-- JEQ @CONFERE_LIMITE_MIN2 	# Se for igual, vai para os as dezenas de minuto
		tmp(171) := JMP  &  R0  &  '0'  &  x"ba";	-- JMP @FIM_CONFERE_LIMITE  	# Caso o contrário já retorna
		tmp(172) := LDA  &  R3  &  '0'  &  x"0d";	-- LDA @13, R3      	#Carrega o valor do limite das dezenas de minuto em R3
		tmp(173) := CEQ  &  R3  &  '0'  &  x"03";	-- CEQ @3, R3     	# Compara com as dezenas de minuto
		tmp(174) := JEQ  &  R0  &  '0'  &  x"b0";	-- JEQ @CONFERE_LIMITE_HORA1 	# Se for igual, vai para as unidades de hora
		tmp(175) := JMP  &  R0  &  '0'  &  x"ba";	-- JMP @FIM_CONFERE_LIMITE   	# Caso o contrário já retorna
		tmp(176) := LDA  &  R0  &  '0'  &  x"0e";	-- LDA @14, R0      	# Carrega o valor do limite das unidades de hora em R0
		tmp(177) := CEQ  &  R0  &  '0'  &  x"04";	-- CEQ @4, R0     	# Compara com as unidades de hora
		tmp(178) := JEQ  &  R0  &  '0'  &  x"b4";	-- JEQ @CONFERE_LIMITE_HORA2 	# Se for igual, vai para as dezenas de hora
		tmp(179) := JMP  &  R0  &  '0'  &  x"ba";	-- JMP @FIM_CONFERE_LIMITE 	# Caso o contrário já retorna
		tmp(180) := LDA  &  R1  &  '0'  &  x"0f";	-- LDA @15, R1      	# Carrega o valor do limite das dezenas de hora em R1
		tmp(181) := CEQ  &  R1  &  '0'  &  x"05";	-- CEQ @5, R1     	# Compara com as dezenas de hora
		tmp(182) := JEQ  &  R0  &  '0'  &  x"b8";	-- JEQ @ATIVA_FLAG_DESPERTADOR 	# Se for igual, vai ativar a flag do despertador
		tmp(183) := JMP  &  R0  &  '0'  &  x"ba";	-- JMP @FIM_CONFERE_LIMITE  	# Caso o contrário já retorna
		tmp(184) := LDA  &  R2  &  '0'  &  x"08";	-- LDA @8, R2      	# Carrega o valor 1
		tmp(185) := STA  &  R2  &  '0'  &  x"06";	-- STA @6, R2      	# Armazena o valor 1 na flag do despertador
		tmp(186) := RET  &  R0  &  '0'  &  x"00";	-- RET
		tmp(187) := STA  &  R0  &  '1'  &  x"fe";	-- STA @510, R0    	# Para limpar a leitura do botão 1
		tmp(188) := STA  &  R3  &  '0'  &  x"06";	-- STA @6, R3      	# Carrega a flag do despertador em R3
		tmp(189) := CEQ  &  R3  &  '0'  &  x"07";	-- CEQ @7, R3      	# Compara a flag do despertador com 0
		tmp(190) := JEQ  &  R0  &  '0'  &  x"c2";	-- JEQ @LIM_UNIDADE 	# Se for 0, então começa a configurar
		tmp(191) := LDA  &  R3  &  '0'  &  x"07";	-- LDA @7, R3      	# Se for 1, tem que voltar para 0
		tmp(192) := STA  &  R3  &  '0'  &  x"06";	-- STA @6, R3      	# Guardo 0 na flag do despertador
		tmp(193) := STA  &  R3  &  '1'  &  x"01";	-- STA @257, R3    	# Guardo 0 no LED8
		tmp(194) := LDA  &  R1  &  '0'  &  x"08";	-- LDA @8, R1      	# Carrega 1 em R1
		tmp(195) := STA  &  R1  &  '1'  &  x"00";	-- STA @256, R1    	# Liga o LED 0 ~ 7 dizendo que está pronto pra ler a chave das unidades de segundo
		tmp(196) := LDA  &  R0  &  '1'  &  x"61";	-- LDA @353, R0    	# Carrega a leitura de KEY1 em R0
		tmp(197) := ANDI  &  R0  &  '0'  &  x"01";	-- ANDI @1, R0     	# Depois de fazer a leitura do botão aplica a máscara
		tmp(198) := CEQ  &  R0  &  '0'  &  x"07";	-- CEQ @7, R0      	# Compara com o valor 0
		tmp(199) := LDA  &  R2  &  '1'  &  x"40";	-- LDA @320, R2    	# Lê as chaves e salva o valor delas no R2
		tmp(200) := JEQ  &  R0  &  '0'  &  x"c2";	-- JEQ @LIM_UNIDADE 	# Caso botão não tenha sido apertado volta novamente para ler KEY1
		tmp(201) := STA  &  R2  &  '0'  &  x"0a";	-- STA @10, R2     	# Guarda o valor limite nas unidades de segundo
		tmp(202) := STA  &  R2  &  '1'  &  x"20";	-- STA @288, R2    	# Guarda o valor das unidades de segundo dos segundos em HEX0
		tmp(203) := STA  &  R0  &  '1'  &  x"fe";	-- STA @510, R0    	# Para limpar a leitura do botão 1
		tmp(204) := LDI  &  R1  &  '0'  &  x"02";	-- LDI $2, R1      	# Carrega 2 em R1
		tmp(205) := STA  &  R1  &  '1'  &  x"00";	-- STA @256, R1    	# Liga o LED 0 ~ 7 dizendo que está pronto pra ler a chave das dezenas
		tmp(206) := LDA  &  R0  &  '1'  &  x"61";	-- LDA @353, R0    	# Guarda a leitura de KEY1 em R0
		tmp(207) := ANDI  &  R0  &  '0'  &  x"01";	-- ANDI @1, R0     	# Depois de fazer a leitura do botão aplica a máscara
		tmp(208) := CEQ  &  R0  &  '0'  &  x"07";	-- CEQ @7, R0      	#Compara com o valor 0
		tmp(209) := LDA  &  R2  &  '1'  &  x"40";	-- LDA @320, R2    	# Lê de novo o valor das chaves e salva no R2
		tmp(210) := JEQ  &  R0  &  '0'  &  x"cc";	-- JEQ @LIM_DEZENA 	# Caso botão não tenha sido apertado volta novamente para ler KEY1
		tmp(211) := STA  &  R2  &  '0'  &  x"0b";	-- STA @11, R2     	# Guarda o valor limite nas dezenas
		tmp(212) := STA  &  R2  &  '1'  &  x"21";	-- STA @289, R2    	# Guarda o valor das dezenas dos segundos em HEX1
		tmp(213) := STA  &  R0  &  '1'  &  x"fe";	-- STA @510, R0    	# Para limpar a leitura do botão 1
		tmp(214) := LDI  &  R1  &  '0'  &  x"04";	-- LDI $4, R1      	# Carrega 4 em R1
		tmp(215) := STA  &  R1  &  '1'  &  x"00";	-- STA @256, R1    	# Liga o LED 0 ~ 7 dizendo que está pronto pra ler a chave das centenas
		tmp(216) := LDA  &  R0  &  '1'  &  x"61";	-- LDA @353, R0    	# Guarda a leitura de KEY1
		tmp(217) := ANDI  &  R0  &  '0'  &  x"01";	-- ANDI @1, R0     	# Depois de fazer a leitura do botão aplica a máscara
		tmp(218) := CEQ  &  R0  &  '0'  &  x"07";	-- CEQ @7, R0      	# Compara com o valor 0
		tmp(219) := LDA  &  R2  &  '1'  &  x"40";	-- LDA @320, R2    	# Lê de novo o valor das chaves e salva no R2
		tmp(220) := JEQ  &  R0  &  '0'  &  x"d6";	-- JEQ @LIM_CENTENA  	# Caso botão não tenha sido apertado volta novamente para ler KEY1
		tmp(221) := STA  &  R2  &  '0'  &  x"0c";	-- STA @12, R2     	# Guarda o valor limite nas centenas
		tmp(222) := STA  &  R2  &  '1'  &  x"22";	-- STA @290, R2    	# Guarda o valor das unidades de segundo dos minutos em HEX2
		tmp(223) := STA  &  R0  &  '1'  &  x"fe";	-- STA @510, R0    	# Para limpar a leitura do botão 1
		tmp(224) := LDI  &  R1  &  '0'  &  x"08";	-- LDI $8, R1      	# Carrega 8 em R1
		tmp(225) := STA  &  R1  &  '1'  &  x"00";	-- STA @256, R1    	# Liga o LED 0 ~ 7 dizendo que está pronto pra ler a chave do milhar
		tmp(226) := LDA  &  R0  &  '1'  &  x"61";	-- LDA @353, R0    	# Guarda a leitura de KEY1
		tmp(227) := ANDI  &  R0  &  '0'  &  x"01";	-- ANDI @1, R0     	# Depois de fazer a leitura do botão aplica a máscara
		tmp(228) := CEQ  &  R0  &  '0'  &  x"07";	-- CEQ @7, R0      	# Compara com o valor 0
		tmp(229) := LDA  &  R2  &  '1'  &  x"40";	-- LDA @320, R2    	# Lê de novo o valor das chaves e salva no R2
		tmp(230) := JEQ  &  R0  &  '0'  &  x"e0";	-- JEQ @LIM_MILHAR  	# Caso botão não tenha sido apertado volta novamente para ler KEY1
		tmp(231) := STA  &  R2  &  '0'  &  x"0d";	-- STA @13, R2     	# Guarda o valor limite nos milhares
		tmp(232) := STA  &  R2  &  '1'  &  x"23";	-- STA @291, R2    	# Guarda o valor das dezenas dos minutos em HEX3
		tmp(233) := STA  &  R0  &  '1'  &  x"fe";	-- STA @510, R0    	# Para limpar a leitura do botão 1 
		tmp(234) := LDI  &  R1  &  '0'  &  x"10";	-- LDI $16, R1     	# Carrega 16 em R1
		tmp(235) := STA  &  R1  &  '1'  &  x"00";	-- STA @256, R1    	# Liga o LED 0 ~ 7 dizendo que está pronto pra ler a chave das dezenas de milhar
		tmp(236) := LDA  &  R0  &  '1'  &  x"61";	-- LDA @353, R0    	# Guarda a leitura de KEY1
		tmp(237) := ANDI  &  R0  &  '0'  &  x"01";	-- ANDI @1, R0     	# Depois de fazer a leitura do botão aplica a máscara
		tmp(238) := CEQ  &  R0  &  '0'  &  x"07";	-- CEQ @7, R0      	# Compara com o valor 0
		tmp(239) := LDA  &  R2  &  '1'  &  x"40";	-- LDA @320, R2    	# Lê de novo o valor das chaves e salva no R2
		tmp(240) := JEQ  &  R0  &  '0'  &  x"ea";	-- JEQ @LIM_DEZMILHAR 	# Caso botão não tenha sido apertado volta novamente para ler KEY1
		tmp(241) := STA  &  R2  &  '0'  &  x"0e";	-- STA @14, R2     	# Guarda o valor limite nas dezenas de milhar
		tmp(242) := STA  &  R2  &  '1'  &  x"24";	-- STA @292, R2    	# Guarda o valor das unidades de segundo das horas em HEX4
		tmp(243) := STA  &  R0  &  '1'  &  x"fe";	-- STA @510, R0    	# Para limpar a leitura do botão 1
		tmp(244) := LDI  &  R1  &  '0'  &  x"20";	-- LDI $32, R1     	# Carrega 32 em R0
		tmp(245) := STA  &  R1  &  '1'  &  x"00";	-- STA @256, R1    	# Liga o LED 0 ~ 7 dizendo que está pronto pra ler a chave das unidades de segundo
		tmp(246) := LDA  &  R0  &  '1'  &  x"61";	-- LDA @353, R0    	# Guarda a leitura de KEY1
		tmp(247) := ANDI  &  R0  &  '0'  &  x"01";	-- ANDI @1, R0     	# Depois de fazer a leitura do botão aplica a máscara
		tmp(248) := CEQ  &  R0  &  '0'  &  x"07";	-- CEQ @7, R0      	#Compara com o valor 0
		tmp(249) := LDA  &  R2  &  '1'  &  x"40";	-- LDA @320, R2    	# Lê de novo o valor das chaves e salva no R2
		tmp(250) := JEQ  &  R0  &  '0'  &  x"f4";	-- JEQ @LIM_CENTMILHAR 	# Caso botão não tenha sido apertado volta novamente para ler KEY1
		tmp(251) := STA  &  R2  &  '0'  &  x"0f";	-- STA @15, R2     	# Guarda o valor limite nas centenas de milhar
		tmp(252) := STA  &  R2  &  '1'  &  x"25";	-- STA @293, R2    	# Guarda o valor das dezenas das horas em HEX5
		tmp(253) := STA  &  R0  &  '1'  &  x"fe";	-- STA @510, R0    	# Para limpar a leitura do botão 1
		tmp(254) := LDA  &  R3  &  '0'  &  x"07";	-- LDA @7, R3      	# Carrega o 0 em R3
		tmp(255) := STA  &  R3  &  '1'  &  x"00";	-- STA @256, R3    	# Desliga os LEDS
		tmp(256) := LDA  &  R0  &  '0'  &  x"0e";	-- LDA @14, R0      	# Carrega as unidades de hora em R0
		tmp(257) := LDA  &  R1  &  '0'  &  x"0f";	-- LDA @15, R1      	# Carrega as dezenas de hora em R1
		tmp(258) := LDA  &  R2  &  '0'  &  x"07";	-- LDA @7, R2
		tmp(259) := ADDI  &  R3  &  '0'  &  x"0a";	-- ADDI $10, R3    	# Soma 10 em R3
		tmp(260) := SUBI  &  R1  &  '0'  &  x"01";	-- SUBI $1, R1     	# Subtrai um de R1
		tmp(261) := CEQ  &  R1  &  '0'  &  x"07";	-- CEQ @7, R1     	# Compara 0 com R1
		tmp(262) := JEQ  &  R0  &  '1'  &  x"08";	-- JEQ @CONTINUA_COMPARACAO_LIMITE
		tmp(263) := JMP  &  R0  &  '1'  &  x"03";	-- JMP @LOOP_PARA_CONCAT_HORA_LIMITE
		tmp(264) := SOMA  &  R3  &  '0'  &  x"0e";	-- SOMA @14, R3    	# Soma as unidades de hora com as dezenas de hora
		tmp(265) := CLT  &  R3  &  '0'  &  x"13";	-- CLT @19, R3     	# R3 é menor que 24?
		tmp(266) := JLT  &  R0  &  '1'  &  x"25";	-- JLT @FIM_LIMITE_DESPERTA  	# Se for menor show de bola
		tmp(267) := CEQ  &  R3  &  '0'  &  x"13";	-- CEQ @19, R3     	# Confere se é igual a 24h
		tmp(268) := JEQ  &  R0  &  '1'  &  x"10";	-- JEQ @EH_24_HORAS_LIMITE
		tmp(269) := LDA  &  R0  &  '0'  &  x"08";	-- LDA @8, R0      	# Se não for menor, carrega 1 em R0
		tmp(270) := STA  &  R0  &  '1'  &  x"02";	-- STA @258, R0    	# Acende o LEDR9
		tmp(271) := JMP  &  R0  &  '0'  &  x"c2";	-- JMP @LIM_UNIDADE 	# Vai configurar a hora de novo
		tmp(272) := LDA  &  R0  &  '0'  &  x"08";	-- LDA @8, R0      	# carrega 1 em R0
		tmp(273) := STA  &  R0  &  '1'  &  x"02";	-- STA @258, R0    	# Acende o LEDR9
		tmp(274) := LDA  &  R0  &  '0'  &  x"07";	-- LDA @7, R0      	# Carrega 0 em R0
		tmp(275) := STA  &  R0  &  '0'  &  x"0e";	-- STA @14, R0      	# Seta as unidades de hora para 0
		tmp(276) := STA  &  R0  &  '0'  &  x"0f";	-- STA @15, R0      	# Seta as dezenas de hora para 0
		tmp(277) := LDA  &  R0  &  '0'  &  x"0a";	-- LDA @10, R0      	# Começa a conferir minutos e segundos
		tmp(278) := CEQ  &  R0  &  '0'  &  x"07";	-- CEQ @7, R0      	# Compara com 0, se não for já volta
		tmp(279) := JEQ  &  R0  &  '1'  &  x"19";	-- JEQ @CONFERE_SEG2_LIMITE 
		tmp(280) := JMP  &  R0  &  '0'  &  x"c2";	-- JMP @LIM_UNIDADE
		tmp(281) := LDA  &  R0  &  '0'  &  x"0b";	-- LDA @11, R0      	# Começa a conferir minutos e segundos
		tmp(282) := CEQ  &  R0  &  '0'  &  x"07";	-- CEQ @7, R0      	# Compara com 0, se não for já volta
		tmp(283) := JEQ  &  R0  &  '1'  &  x"1d";	-- JEQ @CONFERE_MIN1_LIMITE  
		tmp(284) := JMP  &  R0  &  '0'  &  x"cc";	-- JMP @LIM_DEZENA
		tmp(285) := LDA  &  R0  &  '0'  &  x"0c";	-- LDA @12, R0      	# Começa a conferir minutos e segundos
		tmp(286) := CEQ  &  R0  &  '0'  &  x"07";	-- CEQ @7, R0      	# Compara com 0, se não for já volta
		tmp(287) := JEQ  &  R0  &  '1'  &  x"21";	-- JEQ @CONFERE_MIN2_LIMITE 
		tmp(288) := JMP  &  R0  &  '0'  &  x"d6";	-- JMP @LIM_CENTENA
		tmp(289) := LDA  &  R0  &  '0'  &  x"0d";	-- LDA @13, R0      	# Começa a conferir minutos e segundos
		tmp(290) := CEQ  &  R0  &  '0'  &  x"07";	-- CEQ @7, R0      	# Compara com 0, se não for já volta
		tmp(291) := JEQ  &  R0  &  '1'  &  x"25";	-- JEQ @FIM_LIMITE_DESPERTA  
		tmp(292) := JMP  &  R0  &  '0'  &  x"e0";	-- JMP @LIM_MILHAR
		tmp(293) := LDA  &  R0  &  '0'  &  x"07";	-- LDA @7, R0      	# Se não for menor, carrega 1 em R0
		tmp(294) := STA  &  R0  &  '1'  &  x"02";	-- STA @258, R0    	# Apaga o LEDR9
		tmp(295) := RET  &  R0  &  '0'  &  x"00";	-- RET
		tmp(296) := STA  &  R0  &  '1'  &  x"fd";	-- STA @509, R0    	# Para limpar a leitura do botão 2
		tmp(297) := LDA  &  R0  &  '0'  &  x"07";	-- LDA @7, R0      	# Carrega 0 no R0
		tmp(298) := STA  &  R0  &  '0'  &  x"06";	-- STA @6, R0      	# Volta a flag do despertador para 0
		tmp(299) := STA  &  R0  &  '1'  &  x"01";	-- STA @257, R0    	# Salva 0 no LED8
		tmp(300) := STA  &  R0  &  '1'  &  x"02";	-- STA @258, R0    	# Salva 0 no LED8
		tmp(301) := LDA  &  R2  &  '0'  &  x"10";	-- LDA @16, R2     	# Carrega 6 em R2
		tmp(302) := STA  &  R2  &  '0'  &  x"0a";	-- STA @10, R2     	# Armazena o valor do R2 em MEM[10] (valor do despertador para UNIDADE DE SEGUNDO)
		tmp(303) := STA  &  R2  &  '0'  &  x"0b";	-- STA @11, R2     	# Armazena o valor do R2 em MEM[11] (valor do despertador para DEZENA DE SEGUNDO)
		tmp(304) := STA  &  R2  &  '0'  &  x"0c";	-- STA @12, R2     	# Armazena o valor do R2 em MEM[12] (valor do despertador para UNIDADE DE MINUTO)
		tmp(305) := STA  &  R2  &  '0'  &  x"0d";	-- STA @13, R2     	# Armazena o valor do R2 em MEM[13] (valor do despertador para DEZENA DE MINUTO)
		tmp(306) := STA  &  R2  &  '0'  &  x"0e";	-- STA @14, R2     	# Armazena o valor do R2 em MEM[14] (valor do despertador para UNIDADE DE HORA)
		tmp(307) := STA  &  R2  &  '0'  &  x"0f";	-- STA @15, R2     	# Armazena o valor do R2 em MEM[15] (valor do despertador para DEZENA DE HORA)
		tmp(308) := RET  &  R0  &  '0'  &  x"00";	-- RET
		tmp(309) := STA  &  R0  &  '1'  &  x"fc";	-- STA @508, R0    	# Para limpar a leitura do botão 3
		tmp(310) := LDA  &  R1  &  '0'  &  x"08";	-- LDA @8, R1      	# Carrega 1 em R1
		tmp(311) := STA  &  R1  &  '1'  &  x"00";	-- STA @256, R1    	# Liga o LED 0 ~ 7 dizendo que está pronto pra ler a chave das unidades de segundo
		tmp(312) := LDA  &  R0  &  '1'  &  x"63";	-- LDA @355, R0    	# Guarda a leitura de KEY3 em R0
		tmp(313) := ANDI  &  R0  &  '0'  &  x"01";	-- ANDI @1, R0     	# Depois de fazer a leitura do botão aplica a máscara
		tmp(314) := CEQ  &  R0  &  '0'  &  x"07";	-- CEQ @7, R0      	#Compara com o valor 0
		tmp(315) := LDA  &  R2  &  '1'  &  x"40";	-- LDA @320, R2    	# Lê as chaves e salva o valor delas no R2
		tmp(316) := JEQ  &  R0  &  '1'  &  x"36";	-- JEQ @CONFIG_SEG1 	# Caso botão não tenha sido apertado volta novamente para ler KEY3
		tmp(317) := STA  &  R2  &  '0'  &  x"00";	-- STA @0, R2     	# Guarda o valor nas unidades de segundo
		tmp(318) := STA  &  R2  &  '1'  &  x"20";	-- STA @288, R2    	# Guarda o valor das unidades de segundo dos segundos em HEX0
		tmp(319) := STA  &  R0  &  '1'  &  x"fc";	-- STA @508, R0    	# Para limpar a leitura do botão 3
		tmp(320) := LDI  &  R1  &  '0'  &  x"02";	-- LDI $2, R1      	# Carrega 2 em R1
		tmp(321) := STA  &  R1  &  '1'  &  x"00";	-- STA @256, R1    	# Liga o LED 0 ~ 7 dizendo que está pronto pra ler a chave das dezenas
		tmp(322) := LDA  &  R0  &  '1'  &  x"63";	-- LDA @355, R0    	# Guarda a leitura de KEY3 em R0
		tmp(323) := ANDI  &  R0  &  '0'  &  x"01";	-- ANDI @1, R0     	# Depois de fazer a leitura do botão aplica a máscara
		tmp(324) := CEQ  &  R0  &  '0'  &  x"07";	-- CEQ @7, R0      	#Compara com o valor 0
		tmp(325) := LDA  &  R2  &  '1'  &  x"40";	-- LDA @320, R2    	# Lê de novo o valor das chaves e salva no R2
		tmp(326) := JEQ  &  R0  &  '1'  &  x"40";	-- JEQ @CONFIG_SEG2 	# Caso botão não tenha sido apertado volta novamente para ler KEY3
		tmp(327) := STA  &  R2  &  '0'  &  x"01";	-- STA @1, R2     	# Guarda o valor nas dezenas
		tmp(328) := STA  &  R2  &  '1'  &  x"21";	-- STA @289, R2    	# Guarda o valor das dezenas dos segundos em HEX1
		tmp(329) := STA  &  R0  &  '1'  &  x"fc";	-- STA @508, R0    	# Para limpar a leitura do botão 3
		tmp(330) := LDI  &  R1  &  '0'  &  x"04";	-- LDI $4, R1      	# Carrega 4 em R1
		tmp(331) := STA  &  R1  &  '1'  &  x"00";	-- STA @256, R1    	# Liga o LED 0 ~ 7 dizendo que está pronto pra ler a chave das centenas
		tmp(332) := LDA  &  R0  &  '1'  &  x"63";	-- LDA @355, R0    	# Guarda a leitura de KEY3
		tmp(333) := ANDI  &  R0  &  '0'  &  x"01";	-- ANDI @1, R0     	# Depois de fazer a leitura do botão aplica a máscara
		tmp(334) := CEQ  &  R0  &  '0'  &  x"07";	-- CEQ @7, R0      	# Compara com o valor 0
		tmp(335) := LDA  &  R2  &  '1'  &  x"40";	-- LDA @320, R2    	# Lê de novo o valor das chaves e salva no R2
		tmp(336) := JEQ  &  R0  &  '1'  &  x"4a";	-- JEQ @CONFIG_MIN1  	# Caso botão não tenha sido apertado volta novamente para ler KEY3
		tmp(337) := STA  &  R2  &  '0'  &  x"02";	-- STA @2, R2     	# Guarda o valor nas centenas
		tmp(338) := STA  &  R2  &  '1'  &  x"22";	-- STA @290, R2    	# Guarda o valor das unidades de segundo dos minutos em HEX2
		tmp(339) := STA  &  R0  &  '1'  &  x"fc";	-- STA @508, R0    	# Para limpar a leitura do botão 3
		tmp(340) := LDI  &  R1  &  '0'  &  x"08";	-- LDI $8, R1      	# Carrega 8 em R1
		tmp(341) := STA  &  R1  &  '1'  &  x"00";	-- STA @256, R1    	# Liga o LED 0 ~ 7 dizendo que está pronto pra ler a chave do milhar
		tmp(342) := LDA  &  R0  &  '1'  &  x"63";	-- LDA @355, R0    	# Guarda a leitura de KEY3
		tmp(343) := ANDI  &  R0  &  '0'  &  x"01";	-- ANDI @1, R0     	# Depois de fazer a leitura do botão aplica a máscara
		tmp(344) := CEQ  &  R0  &  '0'  &  x"07";	-- CEQ @7, R0      	# Compara com o valor 0
		tmp(345) := LDA  &  R2  &  '1'  &  x"40";	-- LDA @320, R2    	# Lê de novo o valor das chaves e salva no R2
		tmp(346) := JEQ  &  R0  &  '1'  &  x"54";	-- JEQ @CONFIG_MIN2  	# Caso botão não tenha sido apertado volta novamente para ler KEY3
		tmp(347) := STA  &  R2  &  '0'  &  x"03";	-- STA @3, R2     	# Guarda o valor nos milhares
		tmp(348) := STA  &  R2  &  '1'  &  x"23";	-- STA @291, R2    	# Guarda o valor das dezenas dos minutos em HEX3
		tmp(349) := STA  &  R0  &  '1'  &  x"fc";	-- STA @508, R0    	# Para limpar a leitura do botão 3 
		tmp(350) := LDI  &  R1  &  '0'  &  x"10";	-- LDI $16, R1     	# Carrega 16 em R1
		tmp(351) := STA  &  R1  &  '1'  &  x"00";	-- STA @256, R1    	# Liga o LED 0 ~ 7 dizendo que está pronto pra ler a chave das dezenas de milhar
		tmp(352) := LDA  &  R0  &  '1'  &  x"63";	-- LDA @355, R0    	# Guarda a leitura de KEY3
		tmp(353) := ANDI  &  R0  &  '0'  &  x"01";	-- ANDI @1, R0     	# Depois de fazer a leitura do botão aplica a máscara
		tmp(354) := CEQ  &  R0  &  '0'  &  x"07";	-- CEQ @7, R0      	# Compara com o valor 0
		tmp(355) := LDA  &  R2  &  '1'  &  x"40";	-- LDA @320, R2    	# Lê de novo o valor das chaves e salva no R2
		tmp(356) := JEQ  &  R0  &  '1'  &  x"5e";	-- JEQ @CONFIG_HORA1 	# Caso botão não tenha sido apertado volta novamente para ler KEY3
		tmp(357) := STA  &  R2  &  '0'  &  x"04";	-- STA @4, R2     	# Guarda o valor nas dezenas de milhar
		tmp(358) := STA  &  R2  &  '1'  &  x"24";	-- STA @292, R2    	# Guarda o valor das unidades de segundo das horas em HEX4
		tmp(359) := STA  &  R0  &  '1'  &  x"fc";	-- STA @508, R0    	# Para limpar a leitura do botão 3
		tmp(360) := LDI  &  R1  &  '0'  &  x"20";	-- LDI $32, R1     	# Carrega 32 em R0
		tmp(361) := STA  &  R1  &  '1'  &  x"00";	-- STA @256, R1    	# Liga o LED 0 ~ 7 dizendo que está pronto pra ler a chave das unidades de segundo
		tmp(362) := LDA  &  R0  &  '1'  &  x"63";	-- LDA @355, R0    	# Guarda a leitura de KEY3
		tmp(363) := ANDI  &  R0  &  '0'  &  x"01";	-- ANDI @1, R0     	# Depois de fazer a leitura do botão aplica a máscara
		tmp(364) := CEQ  &  R0  &  '0'  &  x"07";	-- CEQ @7, R0      	#Compara com o valor 0
		tmp(365) := LDA  &  R2  &  '1'  &  x"40";	-- LDA @320, R2    	# Lê de novo o valor das chaves e salva no R2
		tmp(366) := JEQ  &  R0  &  '1'  &  x"68";	-- JEQ @CONFIG_HORA2 	# Caso botão não tenha sido apertado volta novamente para ler KEY3
		tmp(367) := STA  &  R2  &  '0'  &  x"05";	-- STA @5, R2     	# Guarda o valor nas centenas de milhar
		tmp(368) := STA  &  R2  &  '1'  &  x"25";	-- STA @293, R2    	# Guarda o valor das dezenas das horas em HEX5
		tmp(369) := STA  &  R0  &  '1'  &  x"fc";	-- STA @508, R0    	# Para limpar a leitura do botão 3
		tmp(370) := LDA  &  R3  &  '0'  &  x"07";	-- LDA @7, R3      	# Carrega o 0 em R3
		tmp(371) := STA  &  R3  &  '1'  &  x"00";	-- STA @256, R3    	# Desliga os LEDS
		tmp(372) := LDA  &  R0  &  '0'  &  x"04";	-- LDA @4, R0      	# Carrega as unidades de hora em R0
		tmp(373) := LDA  &  R1  &  '0'  &  x"05";	-- LDA @5, R1      	# Carrega as dezenas de hora em R1
		tmp(374) := LDA  &  R2  &  '0'  &  x"07";	-- LDA @7, R2
		tmp(375) := ADDI  &  R3  &  '0'  &  x"0a";	-- ADDI $10, R3    	# Soma 10 em R3
		tmp(376) := SUBI  &  R1  &  '0'  &  x"01";	-- SUBI $1, R1     	# Subtrai um de R1
		tmp(377) := CEQ  &  R1  &  '0'  &  x"07";	-- CEQ @7, R1     	# Compara 0 com R1
		tmp(378) := JEQ  &  R0  &  '1'  &  x"7c";	-- JEQ @CONTINUA_COMPARACAO
		tmp(379) := JMP  &  R0  &  '1'  &  x"77";	-- JMP @LOOP_PARA_CONCAT_HORA
		tmp(380) := SOMA  &  R3  &  '0'  &  x"04";	-- SOMA @4, R3    	# Soma as unidades de hora com as dezenas de hora
		tmp(381) := CLT  &  R3  &  '0'  &  x"13";	-- CLT @19, R3     	# R3 é menor que 24?
		tmp(382) := JLT  &  R0  &  '1'  &  x"99";	-- JLT @FIM_CONFIG_HORA  	# Se for menor show de bola
		tmp(383) := CEQ  &  R3  &  '0'  &  x"13";	-- CEQ @19, R3     	# Confere se é igual a 24h
		tmp(384) := JEQ  &  R0  &  '1'  &  x"84";	-- JEQ @EH_24_HORAS
		tmp(385) := LDA  &  R0  &  '0'  &  x"08";	-- LDA @8, R0      	# Se não for menor, carrega 1 em R0
		tmp(386) := STA  &  R0  &  '1'  &  x"02";	-- STA @258, R0    	# Acende o LEDR9
		tmp(387) := JMP  &  R0  &  '1'  &  x"5e";	-- JMP @CONFIG_HORA1 	# Vai configurar a hora de novo
		tmp(388) := LDA  &  R0  &  '0'  &  x"08";	-- LDA @8, R0      	# carrega 1 em R0
		tmp(389) := STA  &  R0  &  '1'  &  x"02";	-- STA @258, R0    	# Acende o LEDR9
		tmp(390) := LDA  &  R0  &  '0'  &  x"07";	-- LDA @7, R0      	# Carrega 0 em R0
		tmp(391) := STA  &  R0  &  '0'  &  x"04";	-- STA @4, R0      	# Seta as unidades de hora para 0
		tmp(392) := STA  &  R0  &  '0'  &  x"05";	-- STA @5, R0      	# Seta as dezenas de hora para 0
		tmp(393) := LDA  &  R0  &  '0'  &  x"00";	-- LDA @0, R0      	# Começa a conferir minutos e segundos
		tmp(394) := CEQ  &  R0  &  '0'  &  x"07";	-- CEQ @7, R0      	# Compara com 0, se não for já volta
		tmp(395) := JEQ  &  R0  &  '1'  &  x"8d";	-- JEQ @CONFERE_SEG2 
		tmp(396) := JMP  &  R0  &  '1'  &  x"36";	-- JMP @CONFIG_SEG1
		tmp(397) := LDA  &  R0  &  '0'  &  x"01";	-- LDA @1, R0      	# Começa a conferir minutos e segundos
		tmp(398) := CEQ  &  R0  &  '0'  &  x"07";	-- CEQ @7, R0      	# Compara com 0, se não for já volta
		tmp(399) := JEQ  &  R0  &  '1'  &  x"91";	-- JEQ @CONFERE_MIN1  
		tmp(400) := JMP  &  R0  &  '1'  &  x"40";	-- JMP @CONFIG_SEG2
		tmp(401) := LDA  &  R0  &  '0'  &  x"02";	-- LDA @2, R0      	# Começa a conferir minutos e segundos
		tmp(402) := CEQ  &  R0  &  '0'  &  x"07";	-- CEQ @7, R0      	# Compara com 0, se não for já volta
		tmp(403) := JEQ  &  R0  &  '1'  &  x"95";	-- JEQ @CONFERE_MIN2  
		tmp(404) := JMP  &  R0  &  '1'  &  x"4a";	-- JMP @CONFIG_MIN1
		tmp(405) := LDA  &  R0  &  '0'  &  x"03";	-- LDA @3, R0      	# Começa a conferir minutos e segundos
		tmp(406) := CEQ  &  R0  &  '0'  &  x"07";	-- CEQ @7, R0      	# Compara com 0, se não for já volta
		tmp(407) := JEQ  &  R0  &  '1'  &  x"99";	-- JEQ @FIM_CONFIG_HORA  
		tmp(408) := JMP  &  R0  &  '1'  &  x"54";	-- JMP @CONFIG_MIN2
		tmp(409) := LDA  &  R0  &  '0'  &  x"07";	-- LDA @7, R0      	# Se não for menor, carrega 1 em R0
		tmp(410) := STA  &  R0  &  '1'  &  x"02";	-- STA @258, R0    	# Apaga o LEDR9
		tmp(411) := RET  &  R0  &  '0'  &  x"00";	-- RET





		  return tmp;
		  
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;