LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY DecoderFunct IS
	PORT (
		FUNCT : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		OUTPUT_FUN : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
	);
END ENTITY;


ARCHITECTURE arch_name OF DecoderFunct IS
	CONSTANT ADDR : STD_LOGIC_VECTOR(5 DOWNTO 0) := "100000";
	CONSTANT SUBR : STD_LOGIC_VECTOR(5 DOWNTO 0) := "100010";
	CONSTANT SLT : STD_LOGIC_VECTOR(5 DOWNTO 0) := "101010";
	CONSTANT ANDR : STD_LOGIC_VECTOR(5 DOWNTO 0) := "100100";
	CONSTANT ORR : STD_LOGIC_VECTOR(5 DOWNTO 0) := "100101";
	CONSTANT JR : STD_LOGIC_VECTOR(5 DOWNTO 0) := "001000";

	-- SelMuxJump|SelMuxRtRd|write_REG(1)|habMUX(rt/imediato)|OP(2)|SelMuxMEMULA|habFlagEqual|
	--read_RAM|write_RAM
BEGIN

	OUTPUT_FUN <= "010" WHEN (FUNCT = ADDR) ELSE
		"110" WHEN (FUNCT = SUBR) ELSE
		"000" WHEN (FUNCT = ANDR) ELSE
		"001" WHEN (FUNCT = ORR) ELSE
		"111" WHEN (FUNCT = SLT) ELSE
		"000" WHEN (FUNCT = JR) ELSE
		"010";

END ARCHITECTURE;