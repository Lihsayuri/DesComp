library ieee;
use ieee.std_logic_1164.all;

entity Aula5final is
  -- Total de bits das entradas e saidas
  generic ( larguraDados : natural := 8;
          larguraEnderecos : natural := 8;
        simulacao : boolean := TRUE -- para gravar na placa, altere de TRUE para FALSE
  );
  port   (
    CLOCK_50 : in std_logic;
    KEY: in std_logic_vector(3 downto 0);
    PC_OUT: out std_logic_vector(larguraEnderecos downto 0);
    LEDR  : out std_logic_vector(9 downto 0);
	 REG_OUT: out std_logic_vector(larguraDados-1 downto 0);
	 SEL_MUX_PC : out std_logic_vector (1 downto 0);
	 Palavra : out std_logic_vector(11 downto 0);
	 JMP_FLAG: out std_logic;
	 JEQ_FLAG: out std_logic;
	 JSR_FLAG: out std_logic;
	 RET_FLAG: out std_logic;
	 EQUAL_FLAG: out std_logic
  );
end entity;


architecture arquitetura of Aula5final is

-- Sinais gerais e sinais do PC: 
  signal CLK : std_logic;
  signal proxPC : std_logic_vector (larguraDados downto 0);
  signal saidaSomador : std_logic_vector (larguraDados downto 0);
  signal Endereco : std_logic_vector (larguraDados downto 0);
  signal instruction: std_logic_vector(12 downto 0);
-- opcode(12 downto 9) endereco(8 downto 0) valor(7 downto 0)

-- Sinais do decodificador de instruções para debug
  signal ULA_FLAG : std_logic;
  signal FLAG_EQ : std_logic;
  signal SelMux2: std_logic_vector (1 downto 0);

-- Sinais de saída do MUX, ALU, Memória, Registrador e Decoder 
  signal MUX_OUT: std_logic_vector(larguraDados - 1 downto 0);
  signal REGA_OUT: std_logic_vector(larguraDados - 1 downto 0);
  signal ULA_OUT: std_logic_vector(larguraDados - 1 downto 0);
  signal MEM_OUT: std_logic_vector(larguraDados - 1 downto 0);
  signal decoder_OUT : std_logic_vector(11 downto 0); -- sinais de controle e ler/escrever
  signal saidaRET : std_logic_vector(larguraDados downto 0);

-- Aliases para facilitar a leitura do código: MUX 
  alias MUX_A: std_logic_vector(larguraDados - 1 downto 0) is MEM_OUT; -- MUX0
  alias MUX_B: std_logic_vector(larguraDados - 1 downto 0) is instruction(larguraDados - 1 downto 0); -- MUX1
  alias MUX_PC_0 : std_logic_vector(larguraDados downto 0) is saidaSomador;
  alias MUX_PC_1 : std_logic_vector(larguraDados downto 0) is instruction(8 downto 0);
  alias MUX_PC_2 : std_logic_vector(larguraDados downto 0) is saidaRET;
  alias MUX_PC_3 : std_logic_vector(larguraDados downto 0) is instruction(8 downto 0);

  
  -- Aliases para os sinais de controle: DECODER_OUT
  alias MEM_Write: std_logic is decoder_OUT(0);
  alias MEM_Read: std_logic is decoder_OUT(1);
  alias habFlag: std_logic is decoder_OUT(2);
  alias Operacao_ULA: std_logic_vector(1 downto 0) is decoder_OUT(4 downto 3);
  alias Habilita_A: std_logic is decoder_OUT(5);  
  alias SelMux: std_logic is decoder_OUT(6);
  alias jeq : std_logic is decoder_OUT(7);
  alias jsr : std_logic is decoder_OUT(8);
  alias ret : std_logic is decoder_OUT(9);
  alias jmp: std_logic is decoder_OUT(10);
  alias habEscritaRet: std_logic is decoder_OUT(11);

  
-- Aliases para facilitar a leitura do código: REGA
  alias REGA_IN: std_logic_vector(larguraDados - 1 downto 0) is ULA_OUT;
  
-- Aliases para facilitar a leitura do código: ULA
  alias ULA_A_IN: std_logic_vector(larguraDados - 1 downto 0) is REGA_OUT;
  alias ULA_B_IN: std_logic_vector(larguraDados - 1 downto 0) is MUX_OUT;

-- Aliases para facilitar a leitura do código: Memória
  alias MEM_ADD: std_logic_vector(larguraDados - 1 downto 0) is instruction(larguraDados - 1 downto 0);
  alias MEM_Habilita: std_logic is instruction(8); 
  alias MEM_IN: std_logic_vector(larguraDados - 1 downto 0) is REGA_OUT;  
  alias OP_CODE: std_logic_vector(3 downto 0) is instruction(12 downto 9); 

  
begin


	-- Instanciando os componentes:

	-- Para simular, fica mais simples tirar o edgeDetector
	gravar:  if simulacao generate
	CLK <= KEY(0);
	else generate
	detectorSub0: work.edgeDetector(bordaSubida)
			  port map (
						clk => CLOCK_50,
						entrada => (not KEY(0)),
						saida => CLK);
	end generate;
	
	-- O port map completo do Program Counter.
	PC : entity work.registradorGenerico generic map (larguraDados => larguraEnderecos+1)
				 port map (
							DIN => proxPC,
							DOUT => Endereco,
							ENABLE => '1',
							CLK => CLK,
							RST => '0');

	incrementaPC :  entity work.somaConstante generic map (larguraDados => larguraEnderecos+1, constante => 1)
			  port map( 
						entrada => Endereco,
						saida => saidaSomador);

	REG_RET : entity work.registradorGenerico generic map (larguraDados => larguraDados+1)
				 port map (
						 DIN => saidaSomador,
						 DOUT => saidaRET,
						 ENABLE => habEscritaRet,
						 CLK => CLK,
						 RST => '0');
						
	MUX2 :  entity work.muxGenerico4x1  generic map (larguraDados => larguraDados+1)
	  port map( 
				  E0 => MUX_PC_0,
				  E1 => MUX_PC_1,
				  E2 => MUX_PC_2,
				  E3 => b"0_0000_0000",
				  SEL_MUX => SelMux2,
				  MUX_OUT => proxPC);
				  
	-- Falta acertar o conteudo da ROM (no arquivo memoriaROM.vhd)
	ROM1 : entity work.memoriaROM generic map (dataWidth => 13, addrWidth =>4) -- POR QUE 4?
				 port map (
						 Endereco => Endereco,
						 Dado => instruction);

	-- O port map completo do MUX.
	MUX1 :  entity work.muxGenerico2x1  generic map (larguraDados => larguraDados)
			  port map( 
						  entradaA_MUX => MUX_A,
						  entradaB_MUX =>  MUX_B,
						  seletor_MUX => SelMux,
						  saida_MUX => MUX_OUT);
						  
	-- O port map completo da ULA:
	ULA1 : entity work.ULASomaSub generic map(larguraDados => larguraDados)
				 port map (
						 entradaA => ULA_A_IN,
						 entradaB => ULA_B_IN,
						 saida => ULA_OUT,
						 seletor => Operacao_ULA,
						 flagEqual => ULA_FLAG);	 
						 
	-- O port map completo do Acumulador.
	REGA : entity work.registradorGenerico generic map (larguraDados => larguraDados)
				 port map (
						 DIN => REGA_IN,
						 DOUT => REGA_OUT,
						 ENABLE => Habilita_A,
						 CLK => CLK,
						 RST => '0');
						 
						 
	-- port map do flip flop da flag de comparacao
	FLAG:
		entity work.flipflopGenerico
		port map (
			DIN		=> ULA_FLAG, 
			DOUT		=> FLAG_EQ,
			ENABLE 	=> habFlag,
			CLK 		=> CLK,
			RST 		=> '0'
		);


	LOG_DESVIO: entity work.logica_desvio
						port map(
							JMP => jmp,
							RET => ret,
							JSR => jsr,
							JEQ => jeq,							
							FLAG_EQ => FLAG_EQ,
							SelMuxPC => SelMux2
						);		


	decoderInstru1 : entity work.decoderInstru
			  port map( 
					  opcode => OP_CODE,
					  saida => decoder_OUT);		
					  

						  
	RAM1 : entity work.memoriaRAM generic map (dataWidth => larguraDados, addrWidth => larguraEnderecos)
				 port map (
						 addr => MEM_ADD,
						 we => MEM_Write,
						 re => MEM_Read,
						 habilita => MEM_Habilita,
						 dado_in => MEM_IN,
						 dado_out => MEM_OUT,
						 clk => CLK);				

	PC_OUT <= Endereco (8 downto 0);
	REG_OUT <= REGA_OUT;
	LEDR(larguraDados - 1 downto 0) <= REGA_OUT;
	LEDR(9 downto 8) <= "00";
	SEL_MUX_PC <= SelMux2;
	JMP_FLAG <= jmp;
	JEQ_FLAG <= jeq;
	JSR_FLAG <= jsr;
	RET_FLAG <= ret;	
	EQUAL_FLAG <= FLAG_EQ;	
	Palavra <= decoder_OUT;
	
end architecture;