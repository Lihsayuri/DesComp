library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity meuNome is
	generic (
		dataWidth: natural := 8; -- tamanho do dado (8 bits)     | Declara apenas
		addrWidth: natural := 3 -- tamanho do endereço (entrada) |  os tamanhos
	);
	port (
		-- O fato da interface ser do tipo std_logic auxilia na simulação
		Endereco : in std_logic_vector (addrWidth-1 downto 0); -- Declara as variáveis
		Dado: out std_logic_vector (dataWidth-1 downto 0)
	);
	
end entity;

-- para ler é assíncrona, para escrever é síncrona!
architecture assincrona of meuNome is
	type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);
-- Basicamente dizendo que o bloco de memória é um array com 8 posições e cada 
-- posição com 8 bits

	function initmemory
		-- Inicializa todas as posições da memória com zero:
		return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
	
	begin
		 -- Inicializa os endereços desejados. Os demais endereços conterão o valor zero:
        tmp(0) := x"4C";
        tmp(1) := x"69";
        tmp(2) := x"76";
        tmp(3) := x"69";
        tmp(4) := x"61";
        tmp(5) := x"5F";
        tmp(6) := x"3A";
        tmp(7) := x"29";
        return tmp;
    end initMemory;
	 
	 signal memROM : blocoMemoria := initMemory;
	
	begin
    -- A conversão de tipos para obter o índice do vetor que será acessado:
    Dado <= memROM (to_integer(unsigned(Endereco)));
	 
end architecture;
